

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO pe64_if_else 
  PIN d[63] 
    ANTENNAPARTIALMETALAREA 0.935 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8024 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 1.0618 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5368 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 8.98761 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 46.8914 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via3 ;
    ANTENNAMAXCUTCAR 0.739298 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.7724 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0608 LAYER Metal4 ;
    ANTENNAGATEAREA 0.288 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 11.6696 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 60.9914 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via4 ;
  END d[63]
  PIN d[62] 
    ANTENNAPARTIALMETALAREA 2.521 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9528 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.168 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 16.2676 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 83.5 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[62]
  PIN d[61] 
    ANTENNAPARTIALMETALAREA 1.0632 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4468 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 19 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 98.03 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.572 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.024 LAYER Metal3 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 23.7667 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 123.23 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via3 ;
    ANTENNAMAXCUTCAR 0.816667 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.6506 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4344 LAYER Metal4 ;
    ANTENNAGATEAREA 0.24 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 26.4775 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 137.54 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.816667 LAYER Via4 ;
  END d[61]
  PIN d[60] 
    ANTENNAPARTIALMETALAREA 1.4222 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.308 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 18.6722 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 97.76 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.762222 LAYER Via4 ;
  END d[60]
  PIN d[59] 
    ANTENNAPARTIALMETALAREA 1.941 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9576 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 10.6307 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 54.2737 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.412632 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.6506 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4344 LAYER Metal3 ;
    ANTENNAGATEAREA 0.288 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 12.8897 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 66.1987 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[59]
  PIN d[58] 
    ANTENNAPARTIALMETALAREA 1.5807 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1108 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 10.3387 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 52.3237 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[58]
  PIN d[57] 
    ANTENNAPARTIALMETALAREA 1.138 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8464 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 17.6447 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 94.72 LAYER Metal6 ;
    ANTENNAMAXCUTCAR 1.41556 LAYER Via6 ;
  END d[57]
  PIN d[56] 
    ANTENNAPARTIALMETALAREA 0.6914 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5496 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.0831 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.522 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.7318 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.852 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 10.1523 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 53.7132 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.739298 LAYER Via4 ;
  END d[56]
  PIN d[55] 
    ANTENNAPARTIALMETALAREA 1.5476 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0352 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 17.8767 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 91.66 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.816667 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.2446 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3464 LAYER Metal3 ;
    ANTENNAGATEAREA 0.18 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 19.2356 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 99.14 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.816667 LAYER Via3 ;
  END d[55]
  PIN d[54] 
    ANTENNAPARTIALMETALAREA 1.709 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7768 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 19.2989 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 100.675 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.816667 LAYER Via4 ;
  END d[54]
  PIN d[53] 
    ANTENNAPARTIALMETALAREA 0.8538 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3848 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.0831 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.522 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.4882 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5992 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.288 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 12.6318 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 66.425 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.721389 LAYER Via4 ;
  END d[53]
  PIN d[52] 
    ANTENNAPARTIALMETALAREA 2.126 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9152 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 12.0404 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 61.1737 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[52]
  PIN d[51] 
    ANTENNAPARTIALMETALAREA 1.7886 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2808 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 20.0217 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 103.77 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[51]
  PIN d[50] 
    ANTENNAPARTIALMETALAREA 0.0418 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2088 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 14.5663 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 76.2026 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.66193 LAYER Via5 ;
  END d[50]
  PIN d[49] 
    ANTENNAPARTIALMETALAREA 1.507 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 27.7104 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 143.79 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 1.2648 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5808 LAYER Metal3 ;
    ANTENNAGATEAREA 0.288 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 32.1021 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 166.64 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via3 ;
    ANTENNAMAXCUTCAR 0.721389 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.6912 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER Metal4 ;
    ANTENNAGATEAREA 0.348 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 34.0883 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 177.109 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via4 ;
  END d[49]
  PIN d[48] 
    ANTENNAPARTIALMETALAREA 1.3868 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1136 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 10.65 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 56.01 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[48]
  PIN d[47] 
    ANTENNAPARTIALMETALAREA 1.3842 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1064 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.288 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 12.4215 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 63.7171 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[47]
  PIN d[46] 
    ANTENNAPARTIALMETALAREA 1.4409 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.398 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.24 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 12.3737 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 64.675 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[46]
  PIN d[45] 
    ANTENNAPARTIALMETALAREA 1.0974 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6376 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.288 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 14.4518 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 75.84 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.838056 LAYER Via5 ;
  END d[45]
  PIN d[44] 
    ANTENNAPARTIALMETALAREA 1.138 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8464 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 17.85 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 93.24 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.871111 LAYER Via5 ;
  END d[44]
  PIN d[43] 
    ANTENNAPARTIALMETALAREA 1.7928 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2016 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.288 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 12.2625 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 62.82 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[43]
  PIN d[42] 
    ANTENNAPARTIALMETALAREA 1.138 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8464 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 13.3344 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 68.1 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.435556 LAYER Via3 ;
  END d[42]
  PIN d[41] 
    ANTENNAPARTIALMETALAREA 0.9756 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0112 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.288 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 15.1348 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 79.4825 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.789444 LAYER Via5 ;
  END d[41]
  PIN d[40] 
    ANTENNAPARTIALMETALAREA 1.1786 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0552 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 13.4621 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 68.735 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via3 ;
  END d[40]
  PIN d[39] 
    ANTENNAPARTIALMETALAREA 1.8334 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4104 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 18.1472 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 94.84 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[39]
  PIN d[38] 
    ANTENNAPARTIALMETALAREA 1.9391 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.954 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 13.3403 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 67.8 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[38]
  PIN d[37] 
    ANTENNAPARTIALMETALAREA 1.8432 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4608 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 18.0758 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 92.14 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.49 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.1634 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9288 LAYER Metal3 ;
    ANTENNAGATEAREA 0.18 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 18.9836 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 97.3 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[37]
  PIN d[36] 
    ANTENNAPARTIALMETALAREA 1.0162 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.22 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 15.2142 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 79.55 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via4 ;
  END d[36]
  PIN d[35] 
    ANTENNAPARTIALMETALAREA 1.7193 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.8236 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 13.3817 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 67.67 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[35]
  PIN d[34] 
    ANTENNAPARTIALMETALAREA 1.8334 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4104 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 17.3758 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 88.57 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.49 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.407 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1816 LAYER Metal3 ;
    ANTENNAGATEAREA 0.18 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 19.6369 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 100.69 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[34]
  PIN d[33] 
    ANTENNAPARTIALMETALAREA 0.8132 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.176 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.2481 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3644 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 10.1233 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 55.16 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via3 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.4476 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3904 LAYER Metal4 ;
    ANTENNAGATEAREA 0.18 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 12.61 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 68.44 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via4 ;
  END d[33]
  PIN d[32] 
    ANTENNAPARTIALMETALAREA 1.341 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8904 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 23.6658 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 121.49 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.407 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1816 LAYER Metal3 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 27.0575 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 139.67 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[32]
  PIN d[31] 
    ANTENNAPARTIALMETALAREA 0.7726 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9672 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.0831 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.522 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 1.5844 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2368 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 23.3267 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 123.53 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.816667 LAYER Via4 ;
  END d[31]
  PIN d[30] 
    ANTENNAPARTIALMETALAREA 2.8052 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4144 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 29.27 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 150.82 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[30]
  PIN d[29] 
    ANTENNAPARTIALMETALAREA 1.1665 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9868 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 14.7008 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 74.59 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[29]
  PIN d[28] 
    ANTENNAPARTIALMETALAREA 0.123 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6264 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 24.9617 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 130.99 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 1.14333 LAYER Via4 ;
  END d[28]
  PIN d[27] 
    ANTENNAPARTIALMETALAREA 0.4072 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.088 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 16.3692 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 85.76 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via4 ;
  END d[27]
  PIN d[26] 
    ANTENNAPARTIALMETALAREA 0.2448 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2528 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 17.3367 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 91.39 LAYER Metal6 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via6 ;
  END d[26]
  PIN d[25] 
    ANTENNAPARTIALMETALAREA 1.7496 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9856 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 20.72 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 105.38 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[25]
  PIN d[24] 
    ANTENNAPARTIALMETALAREA 1.6362 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4024 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 14.9508 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 76.67 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[24]
  PIN d[23] 
    ANTENNAPARTIALMETALAREA 1.5564 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 14.34 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 73.85 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[23]
  PIN d[22] 
    ANTENNAPARTIALMETALAREA 1.5466 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9416 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 14.2042 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 72.83 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[22]
  PIN d[21] 
    ANTENNAPARTIALMETALAREA 1.149 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8968 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 13.975 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 70.94 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.326667 LAYER Via2 ;
  END d[21]
  PIN d[20] 
    ANTENNAPARTIALMETALAREA 0.0418 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2088 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 23.6083 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 124.03 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 1.14333 LAYER Via4 ;
  END d[20]
  PIN d[19] 
    ANTENNAPARTIALMETALAREA 1.303 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6888 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 13.6658 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 71.69 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[19]
  PIN d[18] 
    ANTENNAPARTIALMETALAREA 0.0418 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2088 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 16.1825 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 85.47 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via5 ;
  END d[18]
  PIN d[17] 
    ANTENNAPARTIALMETALAREA 1.2218 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2712 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 19.0117 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 99.1 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[17]
  PIN d[16] 
    ANTENNAPARTIALMETALAREA 0.9756 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0112 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 18.1808 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 96.22 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via5 ;
  END d[16]
  PIN d[15] 
    ANTENNAPARTIALMETALAREA 1.2624 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.48 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 13.275 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 69.95 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[15]
  PIN d[14] 
    ANTENNAPARTIALMETALAREA 1.2624 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.48 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 14.1508 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 73.65 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[14]
  PIN d[13] 
    ANTENNAPARTIALMETALAREA 0.7736 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0608 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 22.6775 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 117.82 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.30667 LAYER Via3 ;
  END d[13]
  PIN d[12] 
    ANTENNAPARTIALMETALAREA 1.0162 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.22 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 15.8517 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 83.82 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via5 ;
  END d[12]
  PIN d[11] 
    ANTENNAPARTIALMETALAREA 1.0162 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.22 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 16.375 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 87.83 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via5 ;
  END d[11]
  PIN d[10] 
    ANTENNAPARTIALMETALAREA 1.0162 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.22 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 15.5079 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 82.39 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via5 ;
  END d[10]
  PIN d[9] 
    ANTENNAPARTIALMETALAREA 1.2624 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.48 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 19.5117 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 100.64 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[9]
  PIN d[8] 
    ANTENNAPARTIALMETALAREA 0.8538 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3848 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 15.9292 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 84.65 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via5 ;
  END d[8]
  PIN d[7] 
    ANTENNAPARTIALMETALAREA 1.2608 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5664 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 19.38 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 101.68 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via3 ;
  END d[7]
  PIN d[6] 
    ANTENNAPARTIALMETALAREA 0.935 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8024 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 17.8425 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 94.48 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.98 LAYER Via5 ;
  END d[6]
  PIN d[5] 
    ANTENNAPARTIALMETALAREA 0.4082 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1816 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 23.1258 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 119.53 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.30667 LAYER Via3 ;
  END d[5]
  PIN d[4] 
    ANTENNAPARTIALMETALAREA 0.326 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6704 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 18.725 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 97.42 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.816667 LAYER Via5 ;
  END d[4]
  PIN d[3] 
    ANTENNAPARTIALMETALAREA 0.8944 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5936 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.5881 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1068 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 7.56583 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 41.84 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[3]
  PIN d[2] 
    ANTENNAPARTIALMETALAREA 0.8132 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.176 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 11.9504 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 62.63 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via4 ;
  END d[2]
  PIN d[1] 
    ANTENNAPARTIALMETALAREA 1.2218 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2712 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 21.5571 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 111.22 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER Via2 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via2 ;
    ANTENNAPARTIALMETALAREA 0.3664 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9728 LAYER Metal3 ;
    ANTENNAGATEAREA 0.168 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 23.738 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 122.963 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.653333 LAYER Via3 ;
  END d[1]
  PIN d[0] 
    ANTENNAPARTIALMETALAREA 1.9094 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8136 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 19.1509 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 99.2556 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.362963 LAYER Via3 ;
  END d[0]
  PIN q[5] 
    ANTENNADIFFAREA 0.168 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.544 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9344 LAYER Metal4 ;
  END q[5]
  PIN q[4] 
    ANTENNADIFFAREA 0.1824 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.356 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1104 LAYER Metal3 ;
  END q[4]
  PIN q[3] 
    ANTENNADIFFAREA 0.2976 LAYER Metal2 ; 
    ANTENNAPARTIALMETALAREA 0.9427 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.842 LAYER Metal2 ;
  END q[3]
  PIN q[2] 
    ANTENNADIFFAREA 0.168 LAYER Metal2 ; 
    ANTENNAPARTIALMETALAREA 1.0162 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.22 LAYER Metal2 ;
  END q[2]
  PIN q[1] 
    ANTENNADIFFAREA 0.168 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.2748 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6928 LAYER Metal3 ;
  END q[1]
  PIN q[0] 
    ANTENNADIFFAREA 0.2832 LAYER Metal2 ; 
    ANTENNAPARTIALMETALAREA 1.1478 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8968 LAYER Metal2 ;
  END q[0]
  PIN v 
    ANTENNADIFFAREA 0.2976 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 2.1936 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2752 LAYER Metal5 ;
  END v
END pe64_if_else

END LIBRARY
