/home/install/FOUNDRY/digital/180nm/dig/lef/all.lef