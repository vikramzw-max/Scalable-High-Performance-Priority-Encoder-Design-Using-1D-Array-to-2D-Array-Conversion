

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO pe64_lookahead 
  PIN d[63] 
    ANTENNAPARTIALMETALAREA 4.6984 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.0836 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5189 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 6.82984 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 29.0583 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.59612 LAYER Via34 ;
  END d[63]
  PIN d[62] 
    ANTENNAPARTIALMETALAREA 2.2624 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5648 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 3.5896 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.886 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6203 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 8.54035 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 35.8613 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.411944 LAYER Via34 ;
  END d[62]
  PIN d[61] 
    ANTENNAPARTIALMETALAREA 2.6376 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.282 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6203 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 8.88846 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 37.5455 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.495385 LAYER Via56 ;
  END d[61]
  PIN d[60] 
    ANTENNAPARTIALMETALAREA 1.9544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6956 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 3.00867 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 12.9044 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.104636 LAYER Via34 ;
  END d[60]
  PIN d[59] 
    ANTENNAPARTIALMETALAREA 1.3076 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9502 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 0.2912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3992 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.368 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8328 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5693 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 9.34479 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 39.1112 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.530811 LAYER Via45 ;
  END d[59]
  PIN d[58] 
    ANTENNAPARTIALMETALAREA 5.9808 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6416 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5621 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 7.63748 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 30.1037 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.293645 LAYER Via34 ;
  END d[58]
  PIN d[57] 
    ANTENNAPARTIALMETALAREA 7.2576 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.772 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0187 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 5.60355 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 22.7421 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.126523 LAYER Via34 ;
  END d[57]
  PIN d[56] 
    ANTENNAPARTIALMETALAREA 4.7572 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.0094 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 5.43367 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 22.1705 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0523179 LAYER Via23 ;
  END d[56]
  PIN d[55] 
    ANTENNAPARTIALMETALAREA 3.3376 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6352 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6563 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 4.64303 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 19.4928 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.226426 LAYER Via34 ;
  END d[55]
  PIN d[54] 
    ANTENNAPARTIALMETALAREA 2.996 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.342 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9179 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 4.49948 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 19.5705 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.143269 LAYER Via34 ;
  END d[54]
  PIN d[53] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.95 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5621 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 5.44634 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 23.044 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.380196 LAYER Via56 ;
  END d[53]
  PIN d[52] 
    ANTENNAPARTIALMETALAREA 2.2848 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6496 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 3.2917 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 13.9258 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.104636 LAYER Via34 ;
  END d[52]
  PIN d[51] 
    ANTENNAPARTIALMETALAREA 1.3076 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9502 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5968 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 5.6784 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7936 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5081 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 14.5197 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 59.5094 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.670751 LAYER Via45 ;
  END d[51]
  PIN d[50] 
    ANTENNAPARTIALMETALAREA 1.6212 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1374 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 1.0304 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1976 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.5808 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6384 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6563 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 6.0013 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 26.3294 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.26724 LAYER Via45 ;
  END d[50]
  PIN d[49] 
    ANTENNAPARTIALMETALAREA 2.6152 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1972 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5621 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 4.7639 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 20.5145 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.544016 LAYER Via45 ;
  END d[49]
  PIN d[48] 
    ANTENNAPARTIALMETALAREA 4.784 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.483 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 6.37474 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 28.8376 LAYER Metal6 ;
  END d[48]
  PIN d[47] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6521 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 4.27951 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 18.138 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.375556 LAYER Via34 ;
  END d[47]
  PIN d[46] 
    ANTENNAPARTIALMETALAREA 5.796 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.942 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6521 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 6.3228 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 25.2285 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.228695 LAYER Via34 ;
  END d[46]
  PIN d[45] 
    ANTENNAPARTIALMETALAREA 4.5416 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.49 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0187 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 5.09431 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 22.0187 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.193497 LAYER Via56 ;
  END d[45]
  PIN d[44] 
    ANTENNAPARTIALMETALAREA 2.2848 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6496 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 3.68888 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 15.9972 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.209272 LAYER Via56 ;
  END d[44]
  PIN d[43] 
    ANTENNAPARTIALMETALAREA 5.3704 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3308 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6521 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 7.1126 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 29.531 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.375556 LAYER Via34 ;
  END d[43]
  PIN d[42] 
    ANTENNAPARTIALMETALAREA 3.5308 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3666 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 3.87826 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 15.8003 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAMAXCUTCAR 0.104636 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 1.7696 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.996 LAYER Metal3 ;
    ANTENNAGATEAREA 2.0187 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 4.75486 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 19.2659 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.186072 LAYER Via34 ;
  END d[42]
  PIN d[41] 
    ANTENNAPARTIALMETALAREA 1.9544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6956 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4829 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 5.23329 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 21.6962 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.399884 LAYER Via34 ;
  END d[41]
  PIN d[40] 
    ANTENNAPARTIALMETALAREA 2.576 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.752 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 3.59941 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 15.3204 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.156954 LAYER Via45 ;
  END d[40]
  PIN d[39] 
    ANTENNAPARTIALMETALAREA 4.5556 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2462 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0187 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 3.40607 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 13.9495 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0930361 LAYER Via23 ;
  END d[39]
  PIN d[38] 
    ANTENNAPARTIALMETALAREA 5.3368 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2036 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7411 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 3.17363 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 12.8261 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0523179 LAYER Via23 ;
  END d[38]
  PIN d[37] 
    ANTENNAPARTIALMETALAREA 6.3364 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.9878 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5143 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 3.95099 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 16.3004 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0553101 LAYER Via23 ;
  END d[37]
  PIN d[36] 
    ANTENNAPARTIALMETALAREA 2.59 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.805 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 3.43534 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 14.3483 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0523179 LAYER Via23 ;
  END d[36]
  PIN d[35] 
    ANTENNAPARTIALMETALAREA 6.1236 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.1822 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6515 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 5.06183 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 20.2897 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.188091 LAYER Via23 ;
  END d[35]
  PIN d[34] 
    ANTENNAPARTIALMETALAREA 3.6736 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9072 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6258 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 7.04698 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 27.0336 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAMAXCUTCAR 0.216043 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5968 LAYER Metal3 ;
    ANTENNAGATEAREA 1.9179 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 7.77694 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 29.9517 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.216043 LAYER Via34 ;
  END d[34]
  PIN d[33] 
    ANTENNAPARTIALMETALAREA 4.5696 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2992 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0187 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 3.7047 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 15.2596 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0930361 LAYER Via23 ;
  END d[33]
  PIN d[32] 
    ANTENNAPARTIALMETALAREA 2.4332 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2114 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 3.3242 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 13.8191 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0523179 LAYER Via23 ;
  END d[32]
  PIN d[31] 
    ANTENNAPARTIALMETALAREA 3.948 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.946 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.109 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 4.64862 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 20.7191 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.600614 LAYER Via56 ;
  END d[31]
  PIN d[30] 
    ANTENNAPARTIALMETALAREA 4.4408 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8116 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.857 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 2.93119 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 10.6856 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAMAXCUTCAR 0.0728056 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5968 LAYER Metal3 ;
    ANTENNAGATEAREA 2.2212 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 3.56148 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 14.4964 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.371225 LAYER Via34 ;
  END d[30]
  PIN d[29] 
    ANTENNAPARTIALMETALAREA 5.5552 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0304 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2212 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 6.34682 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 26.8437 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.371225 LAYER Via34 ;
  END d[29]
  PIN d[28] 
    ANTENNAPARTIALMETALAREA 3.3292 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6034 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2164 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 1.95435 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 7.05423 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0304999 LAYER Via23 ;
  END d[28]
  PIN d[27] 
    ANTENNAPARTIALMETALAREA 5.768 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.836 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1594 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 6.79429 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 27.4633 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.44709 LAYER Via34 ;
  END d[27]
  PIN d[26] 
    ANTENNAPARTIALMETALAREA 4.6592 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6384 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5836 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 3.40863 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 13.6088 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.119201 LAYER Via34 ;
  END d[26]
  PIN d[25] 
    ANTENNAPARTIALMETALAREA 5.5552 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0304 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4828 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 5.38101 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 20.9159 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.189704 LAYER Via56 ;
  END d[25]
  PIN d[24] 
    ANTENNAPARTIALMETALAREA 1.7304 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5508 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.857 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 1.95392 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 7.56327 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.145611 LAYER Via56 ;
  END d[24]
  PIN d[23] 
    ANTENNAPARTIALMETALAREA 4.186 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9866 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 8.23212 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 35.5402 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.521605 LAYER Via23 ;
  END d[23]
  PIN d[22] 
    ANTENNAPARTIALMETALAREA 3.6736 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9072 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7285 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 3.53027 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 14.9437 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.288786 LAYER Via45 ;
  END d[22]
  PIN d[21] 
    ANTENNAPARTIALMETALAREA 6.3364 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.9878 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5188 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 4.2129 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 16.7093 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.223545 LAYER Via23 ;
  END d[21]
  PIN d[20] 
    ANTENNAPARTIALMETALAREA 3.514 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.303 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2164 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 2.03773 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 7.36988 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0304999 LAYER Via23 ;
  END d[20]
  PIN d[19] 
    ANTENNAPARTIALMETALAREA 3.346 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.667 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 5.3872 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.988 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2164 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 4.95315 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 20.9719 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.376183 LAYER Via34 ;
  END d[19]
  PIN d[18] 
    ANTENNAPARTIALMETALAREA 3.9872 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.3912 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9179 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 5.21499 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 21.395 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.143269 LAYER Via34 ;
  END d[18]
  PIN d[17] 
    ANTENNAPARTIALMETALAREA 7.3584 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1536 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5549 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 6.81915 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 27.3834 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.25723 LAYER Via23 ;
  END d[17]
  PIN d[16] 
    ANTENNAPARTIALMETALAREA 3.3292 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6034 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.857 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 2.33259 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 8.41949 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.0364028 LAYER Via23 ;
  END d[16]
  PIN d[15] 
    ANTENNAPARTIALMETALAREA 3.5224 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3348 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0122 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 9.81792 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 39.7636 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.385968 LAYER Via56 ;
  END d[15]
  PIN d[14] 
    ANTENNAPARTIALMETALAREA 7.4032 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.0264 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0122 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 11.507 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 45.2971 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.371225 LAYER Via34 ;
  END d[14]
  PIN d[13] 
    ANTENNAPARTIALMETALAREA 2.5088 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7944 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3746 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 7.6264 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 28.8864 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.306998 LAYER Via56 ;
  END d[13]
  PIN d[12] 
    ANTENNAPARTIALMETALAREA 1.7304 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5508 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 11.5292 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 48.5179 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.208642 LAYER Via34 ;
  END d[12]
  PIN d[11] 
    ANTENNAPARTIALMETALAREA 2.9316 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0982 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 0.8456 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.498 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 1.90203 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 8.47842 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAMAXCUTCAR 0.251488 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.8 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8968 LAYER Metal4 ;
    ANTENNAGATEAREA 1.1706 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 5.73927 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 24.5306 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.556837 LAYER Via45 ;
  END d[11]
  PIN d[10] 
    ANTENNAPARTIALMETALAREA 2.4724 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.6566 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.533 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 4.98465 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 21.2319 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.181229 LAYER Via45 ;
  END d[10]
  PIN d[9] 
    ANTENNAPARTIALMETALAREA 4.2364 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3346 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0836 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 7.25086 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 30.467 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.243867 LAYER Via23 ;
  END d[9]
  PIN d[8] 
    ANTENNAPARTIALMETALAREA 4.784 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.483 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 11.4936 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 52.5425 LAYER Metal6 ;
  END d[8]
  PIN d[7] 
    ANTENNAPARTIALMETALAREA 2.4612 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3174 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 1.5568 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1904 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 6.53302 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 27.5796 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAMAXCUTCAR 0.625926 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 3.8976 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.052 LAYER Metal4 ;
    ANTENNAGATEAREA 1.773 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 8.73133 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 36.0692 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.625926 LAYER Via45 ;
  END d[7]
  PIN d[6] 
    ANTENNAPARTIALMETALAREA 2.59 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.805 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 9.47716 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 36.7074 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAMAXCUTCAR 0.417284 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal3 ;
    ANTENNAGATEAREA 0.324 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 9.80556 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 38.8667 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAMAXCUTCAR 0.625926 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 6.9328 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 26.5424 LAYER Metal4 ;
    ANTENNAGATEAREA 0.4536 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 32.5309 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 130.981 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 1.56481 LAYER Via45 ;
  END d[6]
  PIN d[5] 
    ANTENNAPARTIALMETALAREA 8.988 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.026 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9498 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 11.0766 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 43.9548 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.208642 LAYER Via23 ;
  END d[5]
  PIN d[4] 
    ANTENNAPARTIALMETALAREA 2.7468 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3986 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 11.916 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 49.4994 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.625926 LAYER Via45 ;
  END d[4]
  PIN d[3] 
    ANTENNAPARTIALMETALAREA 2.9456 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1512 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 8.80159 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 33.7428 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAMAXCUTCAR 0.335317 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 0.476 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0988 LAYER Metal3 ;
    ANTENNAGATEAREA 0.4032 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 9.98214 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 38.9482 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAMAXCUTCAR 0.502976 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 5.5076 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.147 LAYER Metal4 ;
    ANTENNAGATEAREA 1.0806 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 15.0789 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 58.5178 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.502976 LAYER Via45 ;
  END d[3]
  PIN d[2] 
    ANTENNAPARTIALMETALAREA 8.6044 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.5738 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7056 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 18.8269 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 73.9967 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.670635 LAYER Via45 ;
  END d[2]
  PIN d[1] 
    ANTENNAPARTIALMETALAREA 4.8808 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.7898 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8676 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 13.0609 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 58.2303 LAYER Metal6 ;
  END d[1]
  PIN d[0] 
    ANTENNAPARTIALMETALAREA 2.59 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.805 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 7.60758 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 29.8782 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.167659 LAYER Via23 ;
  END d[0]
  PIN q[5] 
    ANTENNAPARTIALMETALAREA 4.2868 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.2286 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 4.75876 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 19.25 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAMAXCUTCAR 0.104636 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 0.2912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3992 LAYER Metal3 ;
    ANTENNAGATEAREA 1.2921 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 4.98413 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 20.3329 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAMAXCUTCAR 0.156954 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 4.6816 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.02 LAYER Metal4 ;
    ANTENNAGATEAREA 1.9401 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 9.68325 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 39.1825 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.312963 LAYER Via45 ;
  END q[5]
  PIN q[4] 
    ANTENNADIFFAREA 0.5544 LAYER Metal2 ; 
    ANTENNAPARTIALMETALAREA 3.57 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8118 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 8.02454 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 32.1435 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.104321 LAYER Via23 ;
  END q[4]
  PIN q[3] 
    ANTENNAPARTIALMETALAREA 1.9348 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3246 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via23 ;
    ANTENNAPARTIALMETALAREA 10.8248 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2764 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3505 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 7.31494 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 29.1033 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAMAXCUTCAR 0.18526 LAYER Via34 ;
    ANTENNADIFFAREA 2.757 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 10.7744 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.3824 LAYER Metal4 ;
    ANTENNAGATEAREA 3.5256 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 12.3571 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 49.308 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.563333 LAYER Via45 ;
  END q[3]
  PIN q[2] 
    ANTENNADIFFAREA 0.7845 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.7328 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3456 LAYER Metal4 ;
  END q[2]
  PIN q[1] 
    ANTENNADIFFAREA 1.0368 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.8392 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7484 LAYER Metal3 ;
  END q[1]
  PIN q[0] 
    ANTENNADIFFAREA 0.6144 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.7304 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5508 LAYER Metal3 ;
  END q[0]
  PIN v 
    ANTENNADIFFAREA 1.1206 LAYER Metal2 ; 
    ANTENNAPARTIALMETALAREA 3.346 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.667 LAYER Metal2 ;
  END v
END pe64_lookahead

END LIBRARY
