/home/install/FOUNDRY/digital/90nm/dig/lef/gsclib090_translated.lef